----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    21:13:47 04/03/2022 
-- Design Name: 
-- Module Name:    ADDER_INCREMENTOR - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
use ieee.std_logic_signed.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ADDER_INCREMENTOR is

	port( DataInINC: in std_logic_vector(31 downto 0);
		   DataOutINC: out std_logic_vector(31 downto 0));
			
end ADDER_INCREMENTOR;

architecture Behavioral of ADDER_INCREMENTOR is
	
begin

	DataOutINC <= DataInINC + 4;

end Behavioral;

